------------------------------------------------------------
-- School:     University of Massachusetts Dartmouth      --
-- Department: Computer and Electrical Engineering        --
-- Class:      ECE 368 Digital Design                     --
-- Engineer:   Daniel Noyes                               --
--             Massarrah Tannous                          --
------------------------------------------------------------
--
-- Create Date:    Spring 2014
-- Module Name:    UMDRISC_pkg
-- Project Name:   UMD-RISC 24
-- Target Devices: Spartan-3E
-- Tool versions:  Xilinx ISE 14.7
--
-- Description:
--      This package contain's all the constaints for the 
--          RISC architecture
--
-- Notes:
--      [Insert Notes]
--
-- Revision: 
--      0.01  - File Created
--      0.02  - [Insert]
--
-- Additional Comments: 
--      [Insert Comments]
-- 
-----------------------------------------------------------
package UMDRISC_PKG is

	CONSTANT DATA_WIDTH:INTEGER := 24;
	CONSTANT ADDRESS_WIDTH:INTEGER := 10;
	CONSTANT PC_WIDTH:INTEGER := 10;

end UMDRISC_PKG;

package body UMDRISC_PKG is

end UMDRISC_PKG;
